library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
USE ieee.math_real.ALL;

entity I2C_M_S_RX_TB is
end I2C_M_S_RX_TB;

architecture behavior of I2C_M_S_RX_TB is

	constant clk_period	: time := 10 ns;
	constant DATA_WITH	: integer := 8;
	
	-- IC2 MASTER
	
	constant INPUT_CLK_KHZ 			: integer := 50;
	constant BUS_CLK_MHZ 			: integer := 400;
	constant INPUT_CLK_MULTIPLIER : integer := 100;
	constant BUS_CLK_MULTIPLIER 	: integer := 1;
	
	component I2C_M is
		generic (
										--input clock speed from user logic in KHz
			 input_clk				: integer := INPUT_CLK_KHZ;		
										--speed the I2C_M bus (scl) will run at in MHz 
			 bus_clk					: integer := BUS_CLK_MHZ;		   
										--input clock speed from user logic in KHz
			 input_clk_multiplier: integer := INPUT_CLK_MULTIPLIER;			
			 bus_clk_multiplier	: integer := BUS_CLK_MULTIPLIER
		);
		 port(
			 clk       : in     std_logic;                    --system clock
			 reset_n   : in     std_logic;                    --active low reset
			 ena       : in     std_logic;                    --latch in command
			 addr      : in     std_logic_vector(7 downto 0); --address of target slave
			 rw        : in     std_logic;                    --'0' is write, '1' is read
			 data_wr   : in     std_logic_vector(7 downto 0); --data to write to slave
			 reg_rdy	  : out	  std_logic :='0';				  --ready send the register
			 val_rdy	  : out	  std_logic :='0';				  --ready send value of the register
			 busy      : out    std_logic :='0';              --indicates transaction in progress
			 data_rd   : out    std_logic_vector(7 downto 0); --data read from slave
			 ack_error : out 	  std_logic;                    --flag if improper acknowledge from slave
			 sda       : inout  std_logic;                    --serial data output of I2C_M bus
			 scl       : inout  std_logic  --serial clock output of I2C_M bus
		);                   
	end component;

									--system clock
	signal clk_50				: std_logic:= '0';                    
									--active low reset
	signal rst_n				: std_logic:= '0';                  
									--latch in command
	signal i2c_m_ena			: std_logic:= '0';
									--address of target slave
	signal i2c_m_addr_wr		: std_logic_vector(7 downto 0):= (others=> '0'); 
									--'0' is write, '1' is read
	signal i2c_m_rw			: std_logic:= '1';
									--data to write to slave
	signal i2c_m_data_wr		: std_logic_vector(7 downto 0):= (others=> '0'); 
									--ready send the register
	signal i2c_m_reg_rdy				: std_logic :='0';				  
									--ready send value of the register
	signal i2c_m_val_rdy				: std_logic :='0';				  
									--indicates transaction in progress
	signal i2c_m_busy			: std_logic :='0';              
									--data read from slave
	signal i2c_m_data_rd		: std_logic_vector(7 downto 0):= (others => '0');
									--flag if improper acknowledge from slave	
	signal ack_error			: std_logic:= '0';                    
									--serial data output of I2C_M bus
	signal sda					: std_logic:= 'Z'; 
									--serial clock output of I2C_M bus	
	signal scl					: std_logic:= '0';  
			 
	-- I2C SLAVE RX
	
	constant WR 			: std_logic:='0';
								-- 11h (22h) device address
	constant DEVICE	: std_logic_vector(6 downto 0):= "0100011";		
								-- 00h sub address   
	constant ADDR		: std_logic_vector(7 downto 0):= "10111000";	
	constant REGCONF : std_logic_vector(7 downto 0):= "00010011";	
	constant REGRD : std_logic_vector(7 downto 0):= "01110010";	
	signal VALRD : std_logic_vector(7 downto 0);	
			
	component I2C_S_RX is
		generic(
			WR		: std_logic:= WR;
					-- device address
			DADDR	: std_logic_vector(6 downto 0):= DEVICE;		   
					-- sub address
			ADDR	: std_logic_vector(7 downto 0):= ADDR		
		);
		port(
			RST		: in std_logic;
			SCL		: in std_logic;
			SDA		: inout std_logic;
						-- Recepted over i2c data byte
			DOUT		: out std_logic_vector(7 downto 0);			   
			DATA_RDY	: out std_logic 					
		);
	end component;
	  
	signal i2c_s_rx_data			: std_logic_vector(7 downto 0);
	signal i2c_s_rx_data_rdy	: std_logic;								
	
	-- Build an enumerated type for the state machine
	type state_type is (s0, s1, s2, s3, s4, s5);

	-- Register to hold the current state
	signal state : state_type;
		 
	signal data_error: boolean := false;
begin

	-- IC2 MASTER
	
	UUT : I2C_M 	
	port map (	 			 
		clk 			=> clk_50,
		reset_n 		=> rst_n,
		ena 			=> i2c_m_ena,
		addr 			=> i2c_m_addr_wr,
		rw 			=> i2c_m_rw,
		data_wr 		=> i2c_m_data_wr,
		reg_rdy 		=> i2c_m_reg_rdy,
		val_rdy 		=> i2c_m_val_rdy,
		busy 			=> i2c_m_busy,
		data_rd 		=> i2c_m_data_rd,
		ack_error 	=> ack_error,
		sda 			=> sda,
		scl 			=> scl
	); 
	
	-- I2C SLAVE RX
	
	I_I2C_S_RX: I2C_S_RX
	port map (
		SCL 		=> scl,
		RST 		=> rst_n,
		SDA 		=> sda,
		DOUT 		=> i2c_s_rx_data,
		DATA_RDY	=> i2c_s_rx_data_rdy 
	); 	
	
	P_CLK: process 
	begin
		clk_50 <= '1';
		wait for clk_period/2;
		clk_50 <= '0';
		wait for clk_period/2;
	end process;
	
	P_RST_N: process
	begin	
		rst_n <= '0';	
		wait for clk_period*50;
		rst_n <= '1';			
		wait;
	end process;
	 
	P_i2c_m_write : process(rst_n,clk_50)	
	variable data_wr: natural range 0 to 2**DATA_WITH-1;
	begin
		if rst_n = '0' then
			data_error <= false;
			data_wr := 0;
			i2c_m_addr_wr	<= (others => '1');
			i2c_m_data_wr <= (others => '1'); 
			i2c_m_ena <= '0';   
			i2c_m_rw <= '0'; 
		elsif rising_edge(clk_50)then
			case state is
				when s0 => 
					if i2c_m_busy = '0' then    
						state <= s1;           			
						i2c_m_addr_wr <= DEVICE & '0'; 
						i2c_m_rw <= '0';
						--data to be written
						i2c_m_data_wr <= ADDR;
					end if;
				when s1 =>   
					i2c_m_ena <= '1';   
					if i2c_m_reg_rdy = '1' then 
						state <= s2; 
						-- i2c_m_data_wr <= std_logic_vector(to_unsigned(data_wr,DATA_WITH));
						i2c_m_data_wr <= REGCONF;
					end if;
				when s2 => 
					if i2c_m_val_rdy = '1' then    
						i2c_m_ena <= '0';   
						state <= s3;      
					end if;
				when s3 => 
					if i2c_m_busy = '0' then    
						state <= s4;           			
						i2c_m_addr_wr <= DEVICE & '1'; 
						i2c_m_rw <= '1';
						--data to be written
						i2c_m_data_wr <= REGRD;
					end if;
				when s4 =>   
					i2c_m_ena <= '1';   
					if i2c_m_val_rdy = '1' then 
						state <= s5; 
						-- i2c_m_data_wr <= std_logic_vector(to_unsigned(data_wr,DATA_WITH));
						i2c_m_data_wr <= REGRD;
					end if;
				when s5 => 
					if i2c_m_val_rdy = '1' then    
						i2c_m_ena <= '0';  
						VALRD <=i2c_m_data_rd;						
						state <= s3;      
					end if;
				when OTHERS =>  
					state <= s0; 
			end case; 
		end if;
	end process;
	
end behavior;